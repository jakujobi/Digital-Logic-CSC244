module controller(
	input logic CLKb,
	output logic enA, enC, enALU
);

	/*
	* create a sequential controller
	* 	need a counter to keep track of current step (sequential logic!) - always_ff
	*	need a combinational logic circuit to assign outputs based on current step - always_comb
	*/

endmodule 