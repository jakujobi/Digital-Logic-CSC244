// Create an SV file named “seven_seg.sv” that contains one SV module name seven_seg.
// Write structural or behavioral SV to describe the operation of seven segment display driver.
// The description should include at least one “dec416” sub module.
// The module should have 4 input wires and have outputs so that when it is connected to a seven segment display the hex digits 0-F are displayed.

module seven_seg(
    input [3:0] in,
    input enable,        //enable: enable signal
    output logic [15:0] out     //out: 16-bit output signal
);

// wire [3:0] dec_in;
// assign dec_in = (in > 4'd9) ? 4'd15 : in;

// dec416 dec1(.in(dec_in), .out(out));

dec416 decoder (
    .in(in),    //in: 4-bit input signal (connected to in)
    .enable(enable),    //enable: enable signal (connected to enable)
    .out(out)   //out: 16-bit output signal
);


endmodule